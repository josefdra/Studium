library ieee;
use ieee.std_logic_1164.all;

entity MODULE is
    port(x: in  STD_LOGIC_VECTOR(3 downto 0);
         y: in  STD_LOGIC_VECTOR(3 downto 0);         
         sum: out STD_LOGIC_VECTOR(3 downto 0);
         cout: out STD_LOGIC
    );
end MODULE;

architecture STRUCT of MODULE is
--##INSERT YOUR CODE HERE 

--##INSERT YOUR CODE HERE END
end STRUCT;

