library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity module is
  port(a: in STD_LOGIC_VECTOR(3 downto 0);
       shamt: in STD_LOGIC_VECTOR(1 downto 0); --rotamt
       right_rotated: out STD_LOGIC_VECTOR(3 downto 0); 
       left_rotated: out STD_LOGIC_VECTOR(3 downto 0)       
  );
end;

architecture arch of module is
begin
--##INSERT YOUR CODE HERE 

--##INSERT YOUR CODE HERE END
end;
