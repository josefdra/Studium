library ieee;
use ieee.std_logic_1164.all;

entity TB_MODULE is
end TB_MODULE;

architecture TESTBENCH of TB_MODULE is
  constant tbase: time:=10 ns;
  constant tcheck: time:=1 ns;
--##INSERT YOUR CODE HERE

--##INSERT YOUR CODE HERE END
end TESTBENCH;
