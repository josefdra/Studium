library ieee;
use ieee.std_logic_1164.all;

entity MODULE is
  port(a: in  STD_LOGIC_VECTOR(1 downto 0);
       y: out STD_LOGIC_VECTOR(3 downto 0)
  );
end MODULE;

architecture BEHAV of MODULE is
--##INSERT YOUR CODE HERE
begin

   
--##INSERT YOUR CODE HERE END
end BEHAV;

