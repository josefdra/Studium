library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity module is
  port(btn: in std_logic_vector(1 downto 0);
       segments: out std_logic_vector(6 downto 0)     
  );
end;

architecture arch of module is
--##INSERT YOUR CODE HERE 
--##INSERT YOUR CODE HERE END
end;
