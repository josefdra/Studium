library IEEE; 
use IEEE.STD_LOGIC_1164.all;
entity sevenseg is
  port(bin: in  STD_LOGIC_VECTOR(3 downto 0);
    segments: out STD_LOGIC_VECTOR(6 downto 0)
  );
end;

architecture arch of sevenseg is
begin
--##INSERT YOUR CODE HERE 

--##INSERT YOUR CODE HERE END
end;
